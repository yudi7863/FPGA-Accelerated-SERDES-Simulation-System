
module channel (
	clk_clk,
	reset_reset_n,
	channel_module_0_channel_input_signal_in,
	channel_module_0_channel_input_signal_in_valid,
	channel_module_0_channel_output_signal_out,
	channel_module_0_channel_output_signal_out_valid);	

	input		clk_clk;
	input		reset_reset_n;
	input	[7:0]	channel_module_0_channel_input_signal_in;
	input		channel_module_0_channel_input_signal_in_valid;
	output	[7:0]	channel_module_0_channel_output_signal_out;
	output		channel_module_0_channel_output_signal_out_valid;
endmodule
