module rx_standalone_tb ();

endmodule